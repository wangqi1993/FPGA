// Copyright (C) 1991-2012 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 32-bit"
// VERSION		"Version 12.0 Build 178 05/31/2012 SJ Full Version"
// CREATED		"Tue Sep 20 10:09:45 2016"

module hc74154 (
	C,
	G1N,
	G2N,
	A,
	B,
	D,
	O0N,
	O1N,
	O2N,
	O3N,
	O4N,
	O5N,
	O6N,
	O7N,
	O8N,
	O9N,
	O10N,
	O11N,
	O12N,
	O13N,
	O14N,
	O15N
);
input wire	C;
input wire	G1N;
input wire	G2N;
input wire	A;
input wire	B;
input wire	D;
output wire	O0N;
output wire	O1N;
output wire	O2N;
output wire	O3N;
output wire	O4N;
output wire	O5N;
output wire	O6N;
output wire	O7N;
output wire	O8N;
output wire	O9N;
output wire	O10N;
output wire	O11N;
output wire	O12N;
output wire	O13N;
output wire	O14N;
output wire	O15N;

wire	SYNTHESIZED_WIRE_100;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;

assign	SYNTHESIZED_WIRE_103 = 1;



assign	O15N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_105);

assign	O14N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_105);

assign	O13N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_105);

assign	O12N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_105);

assign	O11N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_105);

assign	O10N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_105);

assign	O9N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_105);

assign	O8N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_105);

assign	O7N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_109);

assign	O6N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_109);

assign	O5N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_109);

assign	O4N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_104 & SYNTHESIZED_WIRE_109);

assign	O3N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_109);

assign	O2N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_102 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_109);

assign	O1N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_101 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_109);

assign	O0N = ~(SYNTHESIZED_WIRE_100 & SYNTHESIZED_WIRE_106 & SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_103 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_109);

assign	SYNTHESIZED_WIRE_105 =  ~SYNTHESIZED_WIRE_109;

assign	SYNTHESIZED_WIRE_109 =  ~D;

assign	SYNTHESIZED_WIRE_104 =  ~SYNTHESIZED_WIRE_108;

assign	SYNTHESIZED_WIRE_108 =  ~C;

assign	SYNTHESIZED_WIRE_102 =  ~SYNTHESIZED_WIRE_107;

assign	SYNTHESIZED_WIRE_107 =  ~B;

assign	SYNTHESIZED_WIRE_106 =  ~A;

assign	SYNTHESIZED_WIRE_101 =  ~SYNTHESIZED_WIRE_106;

assign	SYNTHESIZED_WIRE_100 = ~(G1N | G2N);



endmodule
